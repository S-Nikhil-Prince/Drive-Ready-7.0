***PCIe Interview Questions***
------------------------------------------

Difference between PCI & PCI-X
Difference between End Point & Legacy End Point
Define Forward & Backward Compatibility
What is the difference between C/T/S and C/A/B (possibly referring to Control, Timing, and Status / Command, Address, Byte)?
Define PCIe Link & Lane
What does PCIe x8, x16, x32 mean?
Explain about Quality of Service (QoS)
What is the difference between ECRC & LCRC?
What are the responsibilities of LTSSM?
What is PCIe and how is it different from older versions like PCI & PCI-X?
What is the purpose of the Transaction Layer in PCIe?
What is the purpose of the Data Link Layer in PCIe?
What is the difference between TLP & DLLP?
Discuss the Completion Timeout in PCIe.
What is the use of PCIe Configuration Space?
How does PCIe handle Interrupt delivery?
What is the concept of Virtual Channel in PCIe?
Difference between all generations of PCIe.
What is the purpose of the PCIe Root Complex?
Define Upstream & Downstream Port.
What is the concept of ATS (Address Translation Service) in PCIe?