*** AXI Protocol Interview Questions ***
------------------------------------------

1)How handshaking works in AXI protocol?
2)What is narrow transfer in AXI protocol?
3)what is aligned transfer in AXI protocol?
4)What is wrap transaction in AXI protocol?
5)what is meant by decode error in AXI protocol?
6)what are the different types of responses in AXI protocol?
7)what is the difference between out of order and outstanding transaction in AXI protocol?
8)what is slave error in AXI protocol and what are the possible reasons for it?
9)what is date interleaving in AXI protocol?
10)what is deadlock condition in AXI protocol?
11)what is minimu and maximum bus width supported in AXI protocol?
12)why "wdata" is treated as buffered signal in AXI protocol?
13)which channels are exclusive to slave in AXI protocol?
14)In AXI protocol, differentiate between beat/burst/transaction?
15)what is an interconnect and its purpose in AXI protocol?
16)what is lock signal and its uses in AXI protocol?
17)if AXI length is 4, what is the burst length?
18)Differentiate between AXI3 and AXI4?
19)how to ensure data integrity on AXI?
20)what is the use of strobe in AXI?
21)how to terminate a read or write burst in AXI? {Not Possible}
22)can master give last signal in middle of burst
23)list any 5 features of AXI protocol?
24)what is the role of cache memory in AXI protocol?
25)how does axi support retry transaction?