module axi_lite_master(
    
)